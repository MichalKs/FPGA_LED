
//=======================================================
//  Generic binary counter module
//=======================================================

module decoder3x8 (
  sel,
  q
);

//=======================================================
//  PARAMETER declarations
//=======================================================



//=======================================================
//  PORT declarations
//=======================================================

  input   [2:0]         sel;
  output  [7:0]         q;
  
//=======================================================
//  REG/WIRE declarations
//=======================================================  

  wire     [7:0]        q;

//=======================================================
//  Structural coding
//=======================================================  
  
  assign q = ( sel == 3'b000) ? 8'h01:
             ( sel == 3'b001) ? 8'h02:
             ( sel == 3'b010) ? 8'h04:
             ( sel == 3'b011) ? 8'h08:
             ( sel == 3'b100) ? 8'h10:
             ( sel == 3'b101) ? 8'h20:
             ( sel == 3'b110) ? 8'h40:
             8'h80;
             
endmodule
